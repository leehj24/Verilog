library verilog;
use verilog.vl_types.all;
entity lcd_test_vlg_vec_tst is
end lcd_test_vlg_vec_tst;
