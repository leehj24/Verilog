library verilog;
use verilog.vl_types.all;
entity textlcd_vlg_vec_tst is
end textlcd_vlg_vec_tst;
