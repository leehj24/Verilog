library verilog;
use verilog.vl_types.all;
entity mul_vlg_vec_tst is
end mul_vlg_vec_tst;
