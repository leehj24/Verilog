library verilog;
use verilog.vl_types.all;
entity sdiv_vlg_vec_tst is
end sdiv_vlg_vec_tst;
