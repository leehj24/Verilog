module halfadder(sum, cout, a, b);
  output cout, sum;
  input a, b;
  xor(sum,a,b);
  and(cout,a,b);
endmodule
